magic
tech sky130A
magscale 1 2
timestamp 1718312994
<< viali >>
rect 557 765 591 799
rect 833 765 867 799
rect 1109 765 1143 799
rect 1385 765 1419 799
rect 1661 765 1695 799
rect 1937 765 1971 799
rect 2397 765 2431 799
rect 2673 765 2707 799
rect 2949 765 2983 799
rect 3317 765 3351 799
rect 3593 765 3627 799
rect 3869 765 3903 799
rect 4145 765 4179 799
rect 4421 765 4455 799
rect 4789 765 4823 799
rect 5065 765 5099 799
<< metal1 >>
rect 1 2202 5428 2224
rect 1 2150 926 2202
rect 978 2150 990 2202
rect 1042 2150 1054 2202
rect 1106 2150 1118 2202
rect 1170 2150 2326 2202
rect 2378 2150 2390 2202
rect 2442 2150 2454 2202
rect 2506 2150 2518 2202
rect 2570 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 5428 2202
rect 1 2128 5428 2150
rect 1 1658 5428 1680
rect 1 1606 226 1658
rect 278 1606 290 1658
rect 342 1606 354 1658
rect 406 1606 418 1658
rect 470 1606 1626 1658
rect 1678 1606 1690 1658
rect 1742 1606 1754 1658
rect 1806 1606 1818 1658
rect 1870 1606 3026 1658
rect 3078 1606 3090 1658
rect 3142 1606 3154 1658
rect 3206 1606 3218 1658
rect 3270 1606 4426 1658
rect 4478 1606 4490 1658
rect 4542 1606 4554 1658
rect 4606 1606 4618 1658
rect 4670 1606 5428 1658
rect 1 1584 5428 1606
rect 1 1114 5428 1136
rect 1 1062 926 1114
rect 978 1062 990 1114
rect 1042 1062 1054 1114
rect 1106 1062 1118 1114
rect 1170 1062 2326 1114
rect 2378 1062 2390 1114
rect 2442 1062 2454 1114
rect 2506 1062 2518 1114
rect 2570 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 5428 1114
rect 1 1040 5428 1062
rect 407 796 465 805
rect 545 796 603 805
rect 407 768 603 796
rect 407 759 465 768
rect 545 759 603 768
rect 683 796 741 805
rect 821 796 879 805
rect 683 768 879 796
rect 683 759 741 768
rect 821 759 879 768
rect 959 796 1017 805
rect 1097 796 1155 805
rect 959 768 1155 796
rect 959 759 1017 768
rect 1097 759 1155 768
rect 1235 796 1293 805
rect 1373 796 1431 805
rect 1235 768 1431 796
rect 1235 759 1293 768
rect 1373 759 1431 768
rect 1511 796 1569 805
rect 1649 796 1707 805
rect 1511 768 1707 796
rect 1511 759 1569 768
rect 1649 759 1707 768
rect 1787 796 1845 805
rect 1925 796 1983 805
rect 1787 768 1983 796
rect 1787 759 1845 768
rect 1925 759 1983 768
rect 2247 796 2305 805
rect 2385 796 2443 805
rect 2247 768 2443 796
rect 2247 759 2305 768
rect 2385 759 2443 768
rect 2523 796 2581 805
rect 2661 796 2719 805
rect 2523 768 2719 796
rect 2523 759 2581 768
rect 2661 759 2719 768
rect 2799 796 2857 805
rect 2937 796 2995 805
rect 2799 768 2995 796
rect 2799 759 2857 768
rect 2937 759 2995 768
rect 3167 796 3225 805
rect 3305 796 3363 805
rect 3167 768 3363 796
rect 3167 759 3225 768
rect 3305 759 3363 768
rect 3443 796 3501 805
rect 3581 796 3639 805
rect 3443 768 3639 796
rect 3443 759 3501 768
rect 3581 759 3639 768
rect 3719 796 3777 805
rect 3857 796 3915 805
rect 3719 768 3915 796
rect 3719 759 3777 768
rect 3857 759 3915 768
rect 3995 796 4053 805
rect 4133 796 4191 805
rect 3995 768 4191 796
rect 3995 759 4053 768
rect 4133 759 4191 768
rect 4271 796 4329 805
rect 4409 796 4467 805
rect 4271 768 4467 796
rect 4271 759 4329 768
rect 4409 759 4467 768
rect 4639 796 4697 805
rect 4777 796 4835 805
rect 4639 768 4835 796
rect 4639 759 4697 768
rect 4777 759 4835 768
rect 4915 796 4973 805
rect 5053 796 5111 805
rect 4915 768 5111 796
rect 4915 759 4973 768
rect 5053 759 5111 768
rect 563 711 591 759
rect 839 711 867 759
rect 1115 711 1143 759
rect 1391 711 1419 759
rect 1667 711 1695 759
rect 1943 711 1971 759
rect 2403 711 2431 759
rect 2679 711 2707 759
rect 2955 711 2983 759
rect 3319 711 3347 759
rect 3599 711 3627 759
rect 3875 711 3903 759
rect 4151 711 4179 759
rect 4427 711 4455 759
rect 4795 711 4823 759
rect 5071 711 5099 759
rect 554 705 606 711
rect 554 647 606 653
rect 830 705 882 711
rect 830 647 882 653
rect 1106 705 1158 711
rect 1106 647 1158 653
rect 1382 705 1434 711
rect 1382 647 1434 653
rect 1658 705 1710 711
rect 1658 647 1710 653
rect 1934 705 1986 711
rect 1934 647 1986 653
rect 2394 705 2446 711
rect 2394 647 2446 653
rect 2670 705 2722 711
rect 2670 647 2722 653
rect 2946 705 2998 711
rect 2946 647 2998 653
rect 3310 705 3362 711
rect 3310 647 3362 653
rect 3590 705 3642 711
rect 3590 647 3642 653
rect 3866 705 3918 711
rect 3866 647 3918 653
rect 4142 705 4194 711
rect 4142 647 4194 653
rect 4418 705 4470 711
rect 4418 647 4470 653
rect 4786 705 4838 711
rect 4786 647 4838 653
rect 5062 705 5114 711
rect 5062 647 5114 653
rect 1 570 5428 592
rect 1 518 226 570
rect 278 518 290 570
rect 342 518 354 570
rect 406 518 418 570
rect 470 518 1626 570
rect 1678 518 1690 570
rect 1742 518 1754 570
rect 1806 518 1818 570
rect 1870 518 3026 570
rect 3078 518 3090 570
rect 3142 518 3154 570
rect 3206 518 3218 570
rect 3270 518 4426 570
rect 4478 518 4490 570
rect 4542 518 4554 570
rect 4606 518 4618 570
rect 4670 518 5428 570
rect 1 496 5428 518
<< via1 >>
rect 926 2150 978 2202
rect 990 2150 1042 2202
rect 1054 2150 1106 2202
rect 1118 2150 1170 2202
rect 2326 2150 2378 2202
rect 2390 2150 2442 2202
rect 2454 2150 2506 2202
rect 2518 2150 2570 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 226 1606 278 1658
rect 290 1606 342 1658
rect 354 1606 406 1658
rect 418 1606 470 1658
rect 1626 1606 1678 1658
rect 1690 1606 1742 1658
rect 1754 1606 1806 1658
rect 1818 1606 1870 1658
rect 3026 1606 3078 1658
rect 3090 1606 3142 1658
rect 3154 1606 3206 1658
rect 3218 1606 3270 1658
rect 4426 1606 4478 1658
rect 4490 1606 4542 1658
rect 4554 1606 4606 1658
rect 4618 1606 4670 1658
rect 926 1062 978 1114
rect 990 1062 1042 1114
rect 1054 1062 1106 1114
rect 1118 1062 1170 1114
rect 2326 1062 2378 1114
rect 2390 1062 2442 1114
rect 2454 1062 2506 1114
rect 2518 1062 2570 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 554 653 606 705
rect 830 653 882 705
rect 1106 653 1158 705
rect 1382 653 1434 705
rect 1658 653 1710 705
rect 1934 653 1986 705
rect 2394 653 2446 705
rect 2670 653 2722 705
rect 2946 653 2998 705
rect 3310 653 3362 705
rect 3590 653 3642 705
rect 3866 653 3918 705
rect 4142 653 4194 705
rect 4418 653 4470 705
rect 4786 653 4838 705
rect 5062 653 5114 705
rect 226 518 278 570
rect 290 518 342 570
rect 354 518 406 570
rect 418 518 470 570
rect 1626 518 1678 570
rect 1690 518 1742 570
rect 1754 518 1806 570
rect 1818 518 1870 570
rect 3026 518 3078 570
rect 3090 518 3142 570
rect 3154 518 3206 570
rect 3218 518 3270 570
rect 4426 518 4478 570
rect 4490 518 4542 570
rect 4554 518 4606 570
rect 4618 518 4670 570
<< metal2 >>
rect 926 2204 1170 2224
rect 926 2202 940 2204
rect 996 2202 1020 2204
rect 1076 2202 1100 2204
rect 1156 2202 1170 2204
rect 926 2148 940 2150
rect 996 2148 1020 2150
rect 1076 2148 1100 2150
rect 1156 2148 1170 2150
rect 926 2128 1170 2148
rect 2326 2204 2570 2224
rect 2326 2202 2340 2204
rect 2396 2202 2420 2204
rect 2476 2202 2500 2204
rect 2556 2202 2570 2204
rect 2326 2148 2340 2150
rect 2396 2148 2420 2150
rect 2476 2148 2500 2150
rect 2556 2148 2570 2150
rect 2326 2128 2570 2148
rect 3726 2204 3970 2224
rect 3726 2202 3740 2204
rect 3796 2202 3820 2204
rect 3876 2202 3900 2204
rect 3956 2202 3970 2204
rect 3726 2148 3740 2150
rect 3796 2148 3820 2150
rect 3876 2148 3900 2150
rect 3956 2148 3970 2150
rect 3726 2128 3970 2148
rect 226 1660 470 1680
rect 226 1658 240 1660
rect 296 1658 320 1660
rect 376 1658 400 1660
rect 456 1658 470 1660
rect 226 1604 240 1606
rect 296 1604 320 1606
rect 376 1604 400 1606
rect 456 1604 470 1606
rect 226 1584 470 1604
rect 1626 1660 1870 1680
rect 1626 1658 1640 1660
rect 1696 1658 1720 1660
rect 1776 1658 1800 1660
rect 1856 1658 1870 1660
rect 1626 1604 1640 1606
rect 1696 1604 1720 1606
rect 1776 1604 1800 1606
rect 1856 1604 1870 1606
rect 1626 1584 1870 1604
rect 3026 1660 3270 1680
rect 3026 1658 3040 1660
rect 3096 1658 3120 1660
rect 3176 1658 3200 1660
rect 3256 1658 3270 1660
rect 3026 1604 3040 1606
rect 3096 1604 3120 1606
rect 3176 1604 3200 1606
rect 3256 1604 3270 1606
rect 3026 1584 3270 1604
rect 4426 1660 4670 1680
rect 4426 1658 4440 1660
rect 4496 1658 4520 1660
rect 4576 1658 4600 1660
rect 4656 1658 4670 1660
rect 4426 1604 4440 1606
rect 4496 1604 4520 1606
rect 4576 1604 4600 1606
rect 4656 1604 4670 1606
rect 4426 1584 4670 1604
rect 926 1116 1170 1136
rect 926 1114 940 1116
rect 996 1114 1020 1116
rect 1076 1114 1100 1116
rect 1156 1114 1170 1116
rect 926 1060 940 1062
rect 996 1060 1020 1062
rect 1076 1060 1100 1062
rect 1156 1060 1170 1062
rect 926 1040 1170 1060
rect 2326 1116 2570 1136
rect 2326 1114 2340 1116
rect 2396 1114 2420 1116
rect 2476 1114 2500 1116
rect 2556 1114 2570 1116
rect 2326 1060 2340 1062
rect 2396 1060 2420 1062
rect 2476 1060 2500 1062
rect 2556 1060 2570 1062
rect 2326 1040 2570 1060
rect 3726 1116 3970 1136
rect 3726 1114 3740 1116
rect 3796 1114 3820 1116
rect 3876 1114 3900 1116
rect 3956 1114 3970 1116
rect 3726 1060 3740 1062
rect 3796 1060 3820 1062
rect 3876 1060 3900 1062
rect 3956 1060 3970 1062
rect 3726 1040 3970 1060
rect 548 693 554 705
rect 522 653 554 693
rect 606 653 612 705
rect 824 693 830 705
rect 768 665 830 693
rect 226 572 470 592
rect 226 570 240 572
rect 296 570 320 572
rect 376 570 400 572
rect 456 570 470 572
rect 226 516 240 518
rect 296 516 320 518
rect 376 516 400 518
rect 456 516 470 518
rect 226 496 470 516
rect 522 474 550 653
rect 491 445 550 474
rect 491 400 519 445
rect 768 400 796 665
rect 824 653 830 665
rect 882 653 888 705
rect 1100 693 1106 705
rect 1044 665 1106 693
rect 1044 400 1072 665
rect 1100 653 1106 665
rect 1158 653 1164 705
rect 1376 693 1382 705
rect 1320 665 1382 693
rect 1320 400 1348 665
rect 1376 653 1382 665
rect 1434 653 1440 705
rect 1652 693 1658 705
rect 1556 665 1658 693
rect 1556 465 1584 665
rect 1652 653 1658 665
rect 1710 653 1716 705
rect 1928 653 1934 705
rect 1986 653 1992 705
rect 2388 693 2394 705
rect 2332 665 2394 693
rect 1626 572 1870 592
rect 1626 570 1640 572
rect 1696 570 1720 572
rect 1776 570 1800 572
rect 1856 570 1870 572
rect 1626 516 1640 518
rect 1696 516 1720 518
rect 1776 516 1800 518
rect 1856 516 1870 518
rect 1626 496 1870 516
rect 1945 483 1973 653
rect 1556 437 1624 465
rect 1945 453 1992 483
rect 1596 400 1624 437
rect 1964 400 1992 453
rect 2332 400 2360 665
rect 2388 653 2394 665
rect 2446 653 2452 705
rect 2664 693 2670 705
rect 2608 665 2670 693
rect 2608 400 2636 665
rect 2664 653 2670 665
rect 2722 653 2728 705
rect 2940 693 2946 705
rect 2884 665 2946 693
rect 2884 400 2912 665
rect 2940 653 2946 665
rect 2998 653 3004 705
rect 3304 653 3310 705
rect 3362 653 3368 705
rect 3584 693 3590 705
rect 3528 665 3590 693
rect 3026 572 3270 592
rect 3026 570 3040 572
rect 3096 570 3120 572
rect 3176 570 3200 572
rect 3256 570 3270 572
rect 3026 516 3040 518
rect 3096 516 3120 518
rect 3176 516 3200 518
rect 3256 516 3270 518
rect 3026 496 3270 516
rect 3320 459 3348 653
rect 3252 431 3348 459
rect 3252 400 3280 431
rect 3528 400 3556 665
rect 3584 653 3590 665
rect 3642 653 3648 705
rect 3860 693 3866 705
rect 3804 665 3866 693
rect 3804 400 3832 665
rect 3860 653 3866 665
rect 3918 653 3924 705
rect 4136 693 4142 705
rect 4080 665 4142 693
rect 4080 400 4108 665
rect 4136 653 4142 665
rect 4194 653 4200 705
rect 4412 693 4418 705
rect 4356 665 4418 693
rect 4356 400 4384 665
rect 4412 653 4418 665
rect 4470 653 4476 705
rect 4780 693 4786 705
rect 4724 665 4786 693
rect 4426 572 4670 592
rect 4426 570 4440 572
rect 4496 570 4520 572
rect 4576 570 4600 572
rect 4656 570 4670 572
rect 4426 516 4440 518
rect 4496 516 4520 518
rect 4576 516 4600 518
rect 4656 516 4670 518
rect 4426 496 4670 516
rect 4724 400 4752 665
rect 4780 653 4786 665
rect 4838 653 4844 705
rect 5056 693 5062 705
rect 5000 665 5062 693
rect 5000 400 5028 665
rect 5056 653 5062 665
rect 5114 653 5120 705
rect 478 0 534 400
rect 754 0 810 400
rect 1030 0 1086 400
rect 1306 0 1362 400
rect 1582 0 1638 400
rect 1950 0 2006 400
rect 2318 0 2374 400
rect 2594 0 2650 400
rect 2870 0 2926 400
rect 3238 0 3294 400
rect 3514 0 3570 400
rect 3790 0 3846 400
rect 4066 0 4122 400
rect 4342 0 4398 400
rect 4710 0 4766 400
rect 4986 0 5042 400
<< via2 >>
rect 940 2202 996 2204
rect 1020 2202 1076 2204
rect 1100 2202 1156 2204
rect 940 2150 978 2202
rect 978 2150 990 2202
rect 990 2150 996 2202
rect 1020 2150 1042 2202
rect 1042 2150 1054 2202
rect 1054 2150 1076 2202
rect 1100 2150 1106 2202
rect 1106 2150 1118 2202
rect 1118 2150 1156 2202
rect 940 2148 996 2150
rect 1020 2148 1076 2150
rect 1100 2148 1156 2150
rect 2340 2202 2396 2204
rect 2420 2202 2476 2204
rect 2500 2202 2556 2204
rect 2340 2150 2378 2202
rect 2378 2150 2390 2202
rect 2390 2150 2396 2202
rect 2420 2150 2442 2202
rect 2442 2150 2454 2202
rect 2454 2150 2476 2202
rect 2500 2150 2506 2202
rect 2506 2150 2518 2202
rect 2518 2150 2556 2202
rect 2340 2148 2396 2150
rect 2420 2148 2476 2150
rect 2500 2148 2556 2150
rect 3740 2202 3796 2204
rect 3820 2202 3876 2204
rect 3900 2202 3956 2204
rect 3740 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3796 2202
rect 3820 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3876 2202
rect 3900 2150 3906 2202
rect 3906 2150 3918 2202
rect 3918 2150 3956 2202
rect 3740 2148 3796 2150
rect 3820 2148 3876 2150
rect 3900 2148 3956 2150
rect 240 1658 296 1660
rect 320 1658 376 1660
rect 400 1658 456 1660
rect 240 1606 278 1658
rect 278 1606 290 1658
rect 290 1606 296 1658
rect 320 1606 342 1658
rect 342 1606 354 1658
rect 354 1606 376 1658
rect 400 1606 406 1658
rect 406 1606 418 1658
rect 418 1606 456 1658
rect 240 1604 296 1606
rect 320 1604 376 1606
rect 400 1604 456 1606
rect 1640 1658 1696 1660
rect 1720 1658 1776 1660
rect 1800 1658 1856 1660
rect 1640 1606 1678 1658
rect 1678 1606 1690 1658
rect 1690 1606 1696 1658
rect 1720 1606 1742 1658
rect 1742 1606 1754 1658
rect 1754 1606 1776 1658
rect 1800 1606 1806 1658
rect 1806 1606 1818 1658
rect 1818 1606 1856 1658
rect 1640 1604 1696 1606
rect 1720 1604 1776 1606
rect 1800 1604 1856 1606
rect 3040 1658 3096 1660
rect 3120 1658 3176 1660
rect 3200 1658 3256 1660
rect 3040 1606 3078 1658
rect 3078 1606 3090 1658
rect 3090 1606 3096 1658
rect 3120 1606 3142 1658
rect 3142 1606 3154 1658
rect 3154 1606 3176 1658
rect 3200 1606 3206 1658
rect 3206 1606 3218 1658
rect 3218 1606 3256 1658
rect 3040 1604 3096 1606
rect 3120 1604 3176 1606
rect 3200 1604 3256 1606
rect 4440 1658 4496 1660
rect 4520 1658 4576 1660
rect 4600 1658 4656 1660
rect 4440 1606 4478 1658
rect 4478 1606 4490 1658
rect 4490 1606 4496 1658
rect 4520 1606 4542 1658
rect 4542 1606 4554 1658
rect 4554 1606 4576 1658
rect 4600 1606 4606 1658
rect 4606 1606 4618 1658
rect 4618 1606 4656 1658
rect 4440 1604 4496 1606
rect 4520 1604 4576 1606
rect 4600 1604 4656 1606
rect 940 1114 996 1116
rect 1020 1114 1076 1116
rect 1100 1114 1156 1116
rect 940 1062 978 1114
rect 978 1062 990 1114
rect 990 1062 996 1114
rect 1020 1062 1042 1114
rect 1042 1062 1054 1114
rect 1054 1062 1076 1114
rect 1100 1062 1106 1114
rect 1106 1062 1118 1114
rect 1118 1062 1156 1114
rect 940 1060 996 1062
rect 1020 1060 1076 1062
rect 1100 1060 1156 1062
rect 2340 1114 2396 1116
rect 2420 1114 2476 1116
rect 2500 1114 2556 1116
rect 2340 1062 2378 1114
rect 2378 1062 2390 1114
rect 2390 1062 2396 1114
rect 2420 1062 2442 1114
rect 2442 1062 2454 1114
rect 2454 1062 2476 1114
rect 2500 1062 2506 1114
rect 2506 1062 2518 1114
rect 2518 1062 2556 1114
rect 2340 1060 2396 1062
rect 2420 1060 2476 1062
rect 2500 1060 2556 1062
rect 3740 1114 3796 1116
rect 3820 1114 3876 1116
rect 3900 1114 3956 1116
rect 3740 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3796 1114
rect 3820 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3876 1114
rect 3900 1062 3906 1114
rect 3906 1062 3918 1114
rect 3918 1062 3956 1114
rect 3740 1060 3796 1062
rect 3820 1060 3876 1062
rect 3900 1060 3956 1062
rect 240 570 296 572
rect 320 570 376 572
rect 400 570 456 572
rect 240 518 278 570
rect 278 518 290 570
rect 290 518 296 570
rect 320 518 342 570
rect 342 518 354 570
rect 354 518 376 570
rect 400 518 406 570
rect 406 518 418 570
rect 418 518 456 570
rect 240 516 296 518
rect 320 516 376 518
rect 400 516 456 518
rect 1640 570 1696 572
rect 1720 570 1776 572
rect 1800 570 1856 572
rect 1640 518 1678 570
rect 1678 518 1690 570
rect 1690 518 1696 570
rect 1720 518 1742 570
rect 1742 518 1754 570
rect 1754 518 1776 570
rect 1800 518 1806 570
rect 1806 518 1818 570
rect 1818 518 1856 570
rect 1640 516 1696 518
rect 1720 516 1776 518
rect 1800 516 1856 518
rect 3040 570 3096 572
rect 3120 570 3176 572
rect 3200 570 3256 572
rect 3040 518 3078 570
rect 3078 518 3090 570
rect 3090 518 3096 570
rect 3120 518 3142 570
rect 3142 518 3154 570
rect 3154 518 3176 570
rect 3200 518 3206 570
rect 3206 518 3218 570
rect 3218 518 3256 570
rect 3040 516 3096 518
rect 3120 516 3176 518
rect 3200 516 3256 518
rect 4440 570 4496 572
rect 4520 570 4576 572
rect 4600 570 4656 572
rect 4440 518 4478 570
rect 4478 518 4490 570
rect 4490 518 4496 570
rect 4520 518 4542 570
rect 4542 518 4554 570
rect 4554 518 4576 570
rect 4600 518 4606 570
rect 4606 518 4618 570
rect 4618 518 4656 570
rect 4440 516 4496 518
rect 4520 516 4576 518
rect 4600 516 4656 518
<< metal3 >>
rect 908 2208 1188 2209
rect 908 2144 936 2208
rect 1000 2144 1016 2208
rect 1080 2144 1096 2208
rect 1160 2144 1188 2208
rect 908 2143 1188 2144
rect 2308 2208 2588 2209
rect 2308 2144 2336 2208
rect 2400 2144 2416 2208
rect 2480 2144 2496 2208
rect 2560 2144 2588 2208
rect 2308 2143 2588 2144
rect 3708 2208 3988 2209
rect 3708 2144 3736 2208
rect 3800 2144 3816 2208
rect 3880 2144 3896 2208
rect 3960 2144 3988 2208
rect 3708 2143 3988 2144
rect 208 1664 488 1665
rect 208 1600 236 1664
rect 300 1600 316 1664
rect 380 1600 396 1664
rect 460 1600 488 1664
rect 208 1599 488 1600
rect 1608 1664 1888 1665
rect 1608 1600 1636 1664
rect 1700 1600 1716 1664
rect 1780 1600 1796 1664
rect 1860 1600 1888 1664
rect 1608 1599 1888 1600
rect 3008 1664 3288 1665
rect 3008 1600 3036 1664
rect 3100 1600 3116 1664
rect 3180 1600 3196 1664
rect 3260 1600 3288 1664
rect 3008 1599 3288 1600
rect 4408 1664 4688 1665
rect 4408 1600 4436 1664
rect 4500 1600 4516 1664
rect 4580 1600 4596 1664
rect 4660 1600 4688 1664
rect 4408 1599 4688 1600
rect 908 1120 1188 1121
rect 908 1056 936 1120
rect 1000 1056 1016 1120
rect 1080 1056 1096 1120
rect 1160 1056 1188 1120
rect 908 1055 1188 1056
rect 2308 1120 2588 1121
rect 2308 1056 2336 1120
rect 2400 1056 2416 1120
rect 2480 1056 2496 1120
rect 2560 1056 2588 1120
rect 2308 1055 2588 1056
rect 3708 1120 3988 1121
rect 3708 1056 3736 1120
rect 3800 1056 3816 1120
rect 3880 1056 3896 1120
rect 3960 1056 3988 1120
rect 3708 1055 3988 1056
rect 208 576 488 577
rect 208 512 236 576
rect 300 512 316 576
rect 380 512 396 576
rect 460 512 488 576
rect 208 511 488 512
rect 1608 576 1888 577
rect 1608 512 1636 576
rect 1700 512 1716 576
rect 1780 512 1796 576
rect 1860 512 1888 576
rect 1608 511 1888 512
rect 3008 576 3288 577
rect 3008 512 3036 576
rect 3100 512 3116 576
rect 3180 512 3196 576
rect 3260 512 3288 576
rect 3008 511 3288 512
rect 4408 576 4688 577
rect 4408 512 4436 576
rect 4500 512 4516 576
rect 4580 512 4596 576
rect 4660 512 4688 576
rect 4408 511 4688 512
<< via3 >>
rect 936 2204 1000 2208
rect 936 2148 940 2204
rect 940 2148 996 2204
rect 996 2148 1000 2204
rect 936 2144 1000 2148
rect 1016 2204 1080 2208
rect 1016 2148 1020 2204
rect 1020 2148 1076 2204
rect 1076 2148 1080 2204
rect 1016 2144 1080 2148
rect 1096 2204 1160 2208
rect 1096 2148 1100 2204
rect 1100 2148 1156 2204
rect 1156 2148 1160 2204
rect 1096 2144 1160 2148
rect 2336 2204 2400 2208
rect 2336 2148 2340 2204
rect 2340 2148 2396 2204
rect 2396 2148 2400 2204
rect 2336 2144 2400 2148
rect 2416 2204 2480 2208
rect 2416 2148 2420 2204
rect 2420 2148 2476 2204
rect 2476 2148 2480 2204
rect 2416 2144 2480 2148
rect 2496 2204 2560 2208
rect 2496 2148 2500 2204
rect 2500 2148 2556 2204
rect 2556 2148 2560 2204
rect 2496 2144 2560 2148
rect 3736 2204 3800 2208
rect 3736 2148 3740 2204
rect 3740 2148 3796 2204
rect 3796 2148 3800 2204
rect 3736 2144 3800 2148
rect 3816 2204 3880 2208
rect 3816 2148 3820 2204
rect 3820 2148 3876 2204
rect 3876 2148 3880 2204
rect 3816 2144 3880 2148
rect 3896 2204 3960 2208
rect 3896 2148 3900 2204
rect 3900 2148 3956 2204
rect 3956 2148 3960 2204
rect 3896 2144 3960 2148
rect 236 1660 300 1664
rect 236 1604 240 1660
rect 240 1604 296 1660
rect 296 1604 300 1660
rect 236 1600 300 1604
rect 316 1660 380 1664
rect 316 1604 320 1660
rect 320 1604 376 1660
rect 376 1604 380 1660
rect 316 1600 380 1604
rect 396 1660 460 1664
rect 396 1604 400 1660
rect 400 1604 456 1660
rect 456 1604 460 1660
rect 396 1600 460 1604
rect 1636 1660 1700 1664
rect 1636 1604 1640 1660
rect 1640 1604 1696 1660
rect 1696 1604 1700 1660
rect 1636 1600 1700 1604
rect 1716 1660 1780 1664
rect 1716 1604 1720 1660
rect 1720 1604 1776 1660
rect 1776 1604 1780 1660
rect 1716 1600 1780 1604
rect 1796 1660 1860 1664
rect 1796 1604 1800 1660
rect 1800 1604 1856 1660
rect 1856 1604 1860 1660
rect 1796 1600 1860 1604
rect 3036 1660 3100 1664
rect 3036 1604 3040 1660
rect 3040 1604 3096 1660
rect 3096 1604 3100 1660
rect 3036 1600 3100 1604
rect 3116 1660 3180 1664
rect 3116 1604 3120 1660
rect 3120 1604 3176 1660
rect 3176 1604 3180 1660
rect 3116 1600 3180 1604
rect 3196 1660 3260 1664
rect 3196 1604 3200 1660
rect 3200 1604 3256 1660
rect 3256 1604 3260 1660
rect 3196 1600 3260 1604
rect 4436 1660 4500 1664
rect 4436 1604 4440 1660
rect 4440 1604 4496 1660
rect 4496 1604 4500 1660
rect 4436 1600 4500 1604
rect 4516 1660 4580 1664
rect 4516 1604 4520 1660
rect 4520 1604 4576 1660
rect 4576 1604 4580 1660
rect 4516 1600 4580 1604
rect 4596 1660 4660 1664
rect 4596 1604 4600 1660
rect 4600 1604 4656 1660
rect 4656 1604 4660 1660
rect 4596 1600 4660 1604
rect 936 1116 1000 1120
rect 936 1060 940 1116
rect 940 1060 996 1116
rect 996 1060 1000 1116
rect 936 1056 1000 1060
rect 1016 1116 1080 1120
rect 1016 1060 1020 1116
rect 1020 1060 1076 1116
rect 1076 1060 1080 1116
rect 1016 1056 1080 1060
rect 1096 1116 1160 1120
rect 1096 1060 1100 1116
rect 1100 1060 1156 1116
rect 1156 1060 1160 1116
rect 1096 1056 1160 1060
rect 2336 1116 2400 1120
rect 2336 1060 2340 1116
rect 2340 1060 2396 1116
rect 2396 1060 2400 1116
rect 2336 1056 2400 1060
rect 2416 1116 2480 1120
rect 2416 1060 2420 1116
rect 2420 1060 2476 1116
rect 2476 1060 2480 1116
rect 2416 1056 2480 1060
rect 2496 1116 2560 1120
rect 2496 1060 2500 1116
rect 2500 1060 2556 1116
rect 2556 1060 2560 1116
rect 2496 1056 2560 1060
rect 3736 1116 3800 1120
rect 3736 1060 3740 1116
rect 3740 1060 3796 1116
rect 3796 1060 3800 1116
rect 3736 1056 3800 1060
rect 3816 1116 3880 1120
rect 3816 1060 3820 1116
rect 3820 1060 3876 1116
rect 3876 1060 3880 1116
rect 3816 1056 3880 1060
rect 3896 1116 3960 1120
rect 3896 1060 3900 1116
rect 3900 1060 3956 1116
rect 3956 1060 3960 1116
rect 3896 1056 3960 1060
rect 236 572 300 576
rect 236 516 240 572
rect 240 516 296 572
rect 296 516 300 572
rect 236 512 300 516
rect 316 572 380 576
rect 316 516 320 572
rect 320 516 376 572
rect 376 516 380 572
rect 316 512 380 516
rect 396 572 460 576
rect 396 516 400 572
rect 400 516 456 572
rect 456 516 460 572
rect 396 512 460 516
rect 1636 572 1700 576
rect 1636 516 1640 572
rect 1640 516 1696 572
rect 1696 516 1700 572
rect 1636 512 1700 516
rect 1716 572 1780 576
rect 1716 516 1720 572
rect 1720 516 1776 572
rect 1776 516 1780 572
rect 1716 512 1780 516
rect 1796 572 1860 576
rect 1796 516 1800 572
rect 1800 516 1856 572
rect 1856 516 1860 572
rect 1796 512 1860 516
rect 3036 572 3100 576
rect 3036 516 3040 572
rect 3040 516 3096 572
rect 3096 516 3100 572
rect 3036 512 3100 516
rect 3116 572 3180 576
rect 3116 516 3120 572
rect 3120 516 3176 572
rect 3176 516 3180 572
rect 3116 512 3180 516
rect 3196 572 3260 576
rect 3196 516 3200 572
rect 3200 516 3256 572
rect 3256 516 3260 572
rect 3196 512 3260 516
rect 4436 572 4500 576
rect 4436 516 4440 572
rect 4440 516 4496 572
rect 4496 516 4500 572
rect 4436 512 4500 516
rect 4516 572 4580 576
rect 4516 516 4520 572
rect 4520 516 4576 572
rect 4576 516 4580 572
rect 4516 512 4580 516
rect 4596 572 4660 576
rect 4596 516 4600 572
rect 4600 516 4656 572
rect 4656 516 4660 572
rect 4596 512 4660 516
<< metal4 >>
rect 208 1714 488 2224
rect 208 1478 230 1714
rect 466 1478 488 1714
rect 208 576 488 1478
rect 208 512 236 576
rect 300 512 316 576
rect 380 512 396 576
rect 460 512 488 576
rect 208 496 488 512
rect 908 2208 1188 2224
rect 908 2144 936 2208
rect 1000 2144 1016 2208
rect 1080 2144 1096 2208
rect 1160 2144 1188 2208
rect 908 1120 1188 2144
rect 908 1056 936 1120
rect 1000 1056 1016 1120
rect 1080 1056 1096 1120
rect 1160 1056 1188 1120
rect 908 1014 1188 1056
rect 908 778 930 1014
rect 1166 778 1188 1014
rect 908 496 1188 778
rect 1608 1714 1888 2224
rect 1608 1478 1630 1714
rect 1866 1478 1888 1714
rect 1608 576 1888 1478
rect 1608 512 1636 576
rect 1700 512 1716 576
rect 1780 512 1796 576
rect 1860 512 1888 576
rect 1608 496 1888 512
rect 2308 2208 2588 2224
rect 2308 2144 2336 2208
rect 2400 2144 2416 2208
rect 2480 2144 2496 2208
rect 2560 2144 2588 2208
rect 2308 1120 2588 2144
rect 2308 1056 2336 1120
rect 2400 1056 2416 1120
rect 2480 1056 2496 1120
rect 2560 1056 2588 1120
rect 2308 1014 2588 1056
rect 2308 778 2330 1014
rect 2566 778 2588 1014
rect 2308 496 2588 778
rect 3008 1714 3288 2224
rect 3008 1478 3030 1714
rect 3266 1478 3288 1714
rect 3008 576 3288 1478
rect 3008 512 3036 576
rect 3100 512 3116 576
rect 3180 512 3196 576
rect 3260 512 3288 576
rect 3008 496 3288 512
rect 3708 2208 3988 2224
rect 3708 2144 3736 2208
rect 3800 2144 3816 2208
rect 3880 2144 3896 2208
rect 3960 2144 3988 2208
rect 3708 1120 3988 2144
rect 3708 1056 3736 1120
rect 3800 1056 3816 1120
rect 3880 1056 3896 1120
rect 3960 1056 3988 1120
rect 3708 1014 3988 1056
rect 3708 778 3730 1014
rect 3966 778 3988 1014
rect 3708 496 3988 778
rect 4408 1714 4688 2224
rect 4408 1478 4430 1714
rect 4666 1478 4688 1714
rect 4408 576 4688 1478
rect 4408 512 4436 576
rect 4500 512 4516 576
rect 4580 512 4596 576
rect 4660 512 4688 576
rect 4408 496 4688 512
<< via4 >>
rect 230 1664 466 1714
rect 230 1600 236 1664
rect 236 1600 300 1664
rect 300 1600 316 1664
rect 316 1600 380 1664
rect 380 1600 396 1664
rect 396 1600 460 1664
rect 460 1600 466 1664
rect 230 1478 466 1600
rect 930 778 1166 1014
rect 1630 1664 1866 1714
rect 1630 1600 1636 1664
rect 1636 1600 1700 1664
rect 1700 1600 1716 1664
rect 1716 1600 1780 1664
rect 1780 1600 1796 1664
rect 1796 1600 1860 1664
rect 1860 1600 1866 1664
rect 1630 1478 1866 1600
rect 2330 778 2566 1014
rect 3030 1664 3266 1714
rect 3030 1600 3036 1664
rect 3036 1600 3100 1664
rect 3100 1600 3116 1664
rect 3116 1600 3180 1664
rect 3180 1600 3196 1664
rect 3196 1600 3260 1664
rect 3260 1600 3266 1664
rect 3030 1478 3266 1600
rect 3730 778 3966 1014
rect 4430 1664 4666 1714
rect 4430 1600 4436 1664
rect 4436 1600 4500 1664
rect 4500 1600 4516 1664
rect 4516 1600 4580 1664
rect 4580 1600 4596 1664
rect 4596 1600 4660 1664
rect 4660 1600 4666 1664
rect 4430 1478 4666 1600
<< metal5 >>
rect 1 1714 5428 1756
rect 1 1478 230 1714
rect 466 1478 1630 1714
rect 1866 1478 3030 1714
rect 3266 1478 4430 1714
rect 4666 1478 5428 1714
rect 1 1436 5428 1478
rect 1 1014 5428 1056
rect 1 778 930 1014
rect 1166 778 2330 1014
rect 2566 778 3730 1014
rect 3966 778 5428 1014
rect 1 736 5428 778
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 276 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 276 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1715205430
transform 1 0 2116 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48
timestamp 1715205430
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1715205430
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1715205430
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 4140 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1715205430
transform 1 0 4508 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1715205430
transform 1 0 4692 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1715205430
transform 1 0 5060 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1715205430
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1715205430
transform 1 0 1932 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1715205430
transform 1 0 2116 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1715205430
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 4324 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1715205430
transform 1 0 4692 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp 1715205430
transform 1 0 5060 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_default_value[9] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 3128 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value[10]
timestamp 1715205430
transform 1 0 3404 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value[11]
timestamp 1715205430
transform 1 0 3680 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value[13]
timestamp 1715205430
transform 1 0 4232 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value[14]
timestamp 1715205430
transform 1 0 4600 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value[15]
timestamp 1715205430
transform 1 0 4876 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[0\]
timestamp 1715205430
transform 1 0 368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[1\]
timestamp 1715205430
transform 1 0 644 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[2\]
timestamp 1715205430
transform 1 0 920 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[3\]
timestamp 1715205430
transform 1 0 1196 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[4\]
timestamp 1715205430
transform 1 0 1472 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[5\]
timestamp 1715205430
transform 1 0 1748 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[6\]
timestamp 1715205430
transform 1 0 2208 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[7\]
timestamp 1715205430
transform 1 0 2484 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[8\]
timestamp 1715205430
transform 1 0 2760 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[12\]
timestamp 1715205430
transform 1 0 3956 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1715205430
transform 1 0 0 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1715205430
transform -1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1715205430
transform 1 0 0 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1715205430
transform -1 0 5428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1715205430
transform 1 0 0 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1715205430
transform -1 0 5428 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1715205430
transform 1 0 276 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 2024 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_7
timestamp 1715205430
transform -1 0 4600 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_8
timestamp 1715205430
transform 1 0 4600 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_9
timestamp 1715205430
transform 1 0 2024 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_10
timestamp 1715205430
transform 1 0 4600 0 1 1632
box -38 -48 130 592
<< labels >>
rlabel metal5 s 0 1436 5428 1756 6 VGND
port 0 nsew ground input
rlabel metal4 s 208 496 488 2224 6 VGND
port 0 nsew ground input
rlabel metal4 s 1608 496 1888 2224 6 VGND
port 0 nsew ground input
rlabel metal4 s 3008 496 3288 2224 6 VGND
port 0 nsew ground input
rlabel metal4 s 4408 496 4688 2224 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 736 5428 1056 6 VPWR
port 1 nsew power input
rlabel metal4 s 908 496 1188 2224 6 VPWR
port 1 nsew power input
rlabel metal4 s 2308 496 2588 2224 6 VPWR
port 1 nsew power input
rlabel metal4 s 3708 496 3988 2224 6 VPWR
port 1 nsew power input
rlabel metal2 s 1950 0 2006 400 6 gpio_defaults[5]
port 7 nsew signal tristate
rlabel metal2 s 2594 0 2650 400 6 gpio_defaults[7]
port 9 nsew signal tristate
rlabel metal2 s 2318 0 2374 400 6 gpio_defaults[6]
port 8 nsew signal tristate
rlabel metal2 s 1582 0 1638 400 6 gpio_defaults[4]
port 6 nsew signal tristate
rlabel metal2 s 1306 0 1362 400 6 gpio_defaults[3]
port 5 nsew signal tristate
rlabel metal2 s 1030 0 1086 400 6 gpio_defaults[2]
port 4 nsew signal tristate
rlabel metal2 s 754 0 810 400 6 gpio_defaults[1]
port 3 nsew signal tristate
rlabel metal2 s 478 0 534 400 6 gpio_defaults[0]
port 2 nsew signal tristate
rlabel metal2 s 2870 0 2926 400 6 gpio_defaults[8]
port 10 nsew signal tristate
rlabel metal2 s 3238 0 3294 400 6 gpio_defaults[9]
port 11 nsew signal tristate
rlabel metal2 s 3514 0 3570 400 6 gpio_defaults[10]
port 12 nsew signal tristate
rlabel metal2 s 3790 0 3846 400 6 gpio_defaults[11]
port 13 nsew signal tristate
rlabel metal2 s 4066 0 4122 400 6 gpio_defaults[12]
port 14 nsew signal tristate
rlabel metal2 s 4342 0 4398 400 6 gpio_defaults[13]
port 15 nsew signal tristate
rlabel metal2 s 4710 0 4766 400 6 gpio_defaults[14]
port 16 nsew signal tristate
rlabel metal2 s 4986 0 5042 400 6 gpio_defaults[15]
port 17 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 5428 2200
<< end >>
