magic
tech sky130A
magscale 1 2
timestamp 1718313015
<< viali >>
rect 557 765 591 799
rect 833 765 867 799
rect 1109 765 1143 799
rect 1385 765 1419 799
rect 1661 765 1695 799
rect 1937 765 1971 799
rect 2397 765 2431 799
rect 2673 765 2707 799
<< metal1 >>
rect 1 2202 3204 2224
rect 1 2150 926 2202
rect 978 2150 990 2202
rect 1042 2150 1054 2202
rect 1106 2150 1118 2202
rect 1170 2150 2326 2202
rect 2378 2150 2390 2202
rect 2442 2150 2454 2202
rect 2506 2150 2518 2202
rect 2570 2150 3204 2202
rect 1 2128 3204 2150
rect 1 1658 3204 1680
rect 1 1606 226 1658
rect 278 1606 290 1658
rect 342 1606 354 1658
rect 406 1606 418 1658
rect 470 1606 1626 1658
rect 1678 1606 1690 1658
rect 1742 1606 1754 1658
rect 1806 1606 1818 1658
rect 1870 1606 3204 1658
rect 1 1584 3204 1606
rect 1 1114 3204 1136
rect 1 1062 926 1114
rect 978 1062 990 1114
rect 1042 1062 1054 1114
rect 1106 1062 1118 1114
rect 1170 1062 2326 1114
rect 2378 1062 2390 1114
rect 2442 1062 2454 1114
rect 2506 1062 2518 1114
rect 2570 1062 3204 1114
rect 1 1040 3204 1062
rect 407 796 465 805
rect 545 796 603 805
rect 407 768 603 796
rect 407 759 465 768
rect 545 759 603 768
rect 683 796 741 805
rect 821 796 879 805
rect 683 768 879 796
rect 683 759 741 768
rect 821 759 879 768
rect 959 796 1017 805
rect 1097 796 1155 805
rect 959 768 1155 796
rect 959 759 1017 768
rect 1097 759 1155 768
rect 1235 796 1293 805
rect 1373 796 1431 805
rect 1235 768 1431 796
rect 1235 759 1293 768
rect 1373 759 1431 768
rect 1511 796 1569 805
rect 1649 796 1707 805
rect 1511 768 1707 796
rect 1511 759 1569 768
rect 1649 759 1707 768
rect 1787 796 1845 805
rect 1925 796 1983 805
rect 1787 768 1983 796
rect 1787 759 1845 768
rect 1925 759 1983 768
rect 2247 796 2305 805
rect 2385 796 2443 805
rect 2247 768 2443 796
rect 2247 759 2305 768
rect 2385 759 2443 768
rect 2523 796 2581 805
rect 2661 796 2719 805
rect 2523 768 2719 796
rect 2523 759 2581 768
rect 2661 759 2719 768
rect 563 711 591 759
rect 839 711 867 759
rect 1115 711 1143 759
rect 1391 711 1419 759
rect 1667 711 1695 759
rect 1943 711 1971 759
rect 2403 711 2431 759
rect 2679 711 2707 759
rect 554 705 606 711
rect 554 647 606 653
rect 830 705 882 711
rect 830 647 882 653
rect 1106 705 1158 711
rect 1106 647 1158 653
rect 1382 705 1434 711
rect 1382 647 1434 653
rect 1658 705 1710 711
rect 1658 647 1710 653
rect 1934 705 1986 711
rect 1934 647 1986 653
rect 2394 705 2446 711
rect 2394 647 2446 653
rect 2670 705 2722 711
rect 2670 647 2722 653
rect 1 570 3204 592
rect 1 518 226 570
rect 278 518 290 570
rect 342 518 354 570
rect 406 518 418 570
rect 470 518 1626 570
rect 1678 518 1690 570
rect 1742 518 1754 570
rect 1806 518 1818 570
rect 1870 518 3204 570
rect 1 496 3204 518
<< via1 >>
rect 926 2150 978 2202
rect 990 2150 1042 2202
rect 1054 2150 1106 2202
rect 1118 2150 1170 2202
rect 2326 2150 2378 2202
rect 2390 2150 2442 2202
rect 2454 2150 2506 2202
rect 2518 2150 2570 2202
rect 226 1606 278 1658
rect 290 1606 342 1658
rect 354 1606 406 1658
rect 418 1606 470 1658
rect 1626 1606 1678 1658
rect 1690 1606 1742 1658
rect 1754 1606 1806 1658
rect 1818 1606 1870 1658
rect 926 1062 978 1114
rect 990 1062 1042 1114
rect 1054 1062 1106 1114
rect 1118 1062 1170 1114
rect 2326 1062 2378 1114
rect 2390 1062 2442 1114
rect 2454 1062 2506 1114
rect 2518 1062 2570 1114
rect 554 653 606 705
rect 830 653 882 705
rect 1106 653 1158 705
rect 1382 653 1434 705
rect 1658 653 1710 705
rect 1934 653 1986 705
rect 2394 653 2446 705
rect 2670 653 2722 705
rect 226 518 278 570
rect 290 518 342 570
rect 354 518 406 570
rect 418 518 470 570
rect 1626 518 1678 570
rect 1690 518 1742 570
rect 1754 518 1806 570
rect 1818 518 1870 570
<< metal2 >>
rect 926 2204 1170 2224
rect 926 2202 940 2204
rect 996 2202 1020 2204
rect 1076 2202 1100 2204
rect 1156 2202 1170 2204
rect 926 2148 940 2150
rect 996 2148 1020 2150
rect 1076 2148 1100 2150
rect 1156 2148 1170 2150
rect 926 2128 1170 2148
rect 2326 2204 2570 2224
rect 2326 2202 2340 2204
rect 2396 2202 2420 2204
rect 2476 2202 2500 2204
rect 2556 2202 2570 2204
rect 2326 2148 2340 2150
rect 2396 2148 2420 2150
rect 2476 2148 2500 2150
rect 2556 2148 2570 2150
rect 2326 2128 2570 2148
rect 226 1660 470 1680
rect 226 1658 240 1660
rect 296 1658 320 1660
rect 376 1658 400 1660
rect 456 1658 470 1660
rect 226 1604 240 1606
rect 296 1604 320 1606
rect 376 1604 400 1606
rect 456 1604 470 1606
rect 226 1584 470 1604
rect 1626 1660 1870 1680
rect 1626 1658 1640 1660
rect 1696 1658 1720 1660
rect 1776 1658 1800 1660
rect 1856 1658 1870 1660
rect 1626 1604 1640 1606
rect 1696 1604 1720 1606
rect 1776 1604 1800 1606
rect 1856 1604 1870 1606
rect 1626 1584 1870 1604
rect 926 1116 1170 1136
rect 926 1114 940 1116
rect 996 1114 1020 1116
rect 1076 1114 1100 1116
rect 1156 1114 1170 1116
rect 926 1060 940 1062
rect 996 1060 1020 1062
rect 1076 1060 1100 1062
rect 1156 1060 1170 1062
rect 926 1040 1170 1060
rect 2326 1116 2570 1136
rect 2326 1114 2340 1116
rect 2396 1114 2420 1116
rect 2476 1114 2500 1116
rect 2556 1114 2570 1116
rect 2326 1060 2340 1062
rect 2396 1060 2420 1062
rect 2476 1060 2500 1062
rect 2556 1060 2570 1062
rect 2326 1040 2570 1060
rect 548 693 554 705
rect 522 653 554 693
rect 606 653 612 705
rect 824 693 830 705
rect 768 665 830 693
rect 226 572 470 592
rect 226 570 240 572
rect 296 570 320 572
rect 376 570 400 572
rect 456 570 470 572
rect 226 516 240 518
rect 296 516 320 518
rect 376 516 400 518
rect 456 516 470 518
rect 226 496 470 516
rect 522 474 550 653
rect 491 445 550 474
rect 491 400 519 445
rect 768 400 796 665
rect 824 653 830 665
rect 882 653 888 705
rect 1100 693 1106 705
rect 1044 665 1106 693
rect 1044 400 1072 665
rect 1100 653 1106 665
rect 1158 653 1164 705
rect 1376 693 1382 705
rect 1320 665 1382 693
rect 1320 400 1348 665
rect 1376 653 1382 665
rect 1434 653 1440 705
rect 1652 693 1658 705
rect 1556 665 1658 693
rect 1556 465 1584 665
rect 1652 653 1658 665
rect 1710 653 1716 705
rect 1928 653 1934 705
rect 1986 653 1992 705
rect 2388 693 2394 705
rect 2332 665 2394 693
rect 1626 572 1870 592
rect 1626 570 1640 572
rect 1696 570 1720 572
rect 1776 570 1800 572
rect 1856 570 1870 572
rect 1626 516 1640 518
rect 1696 516 1720 518
rect 1776 516 1800 518
rect 1856 516 1870 518
rect 1626 496 1870 516
rect 1945 483 1973 653
rect 1556 437 1624 465
rect 1945 453 1992 483
rect 1596 400 1624 437
rect 1964 400 1992 453
rect 2332 400 2360 665
rect 2388 653 2394 665
rect 2446 653 2452 705
rect 2664 693 2670 705
rect 2608 665 2670 693
rect 2608 400 2636 665
rect 2664 653 2670 665
rect 2722 653 2728 705
rect 478 0 534 400
rect 754 0 810 400
rect 1030 0 1086 400
rect 1306 0 1362 400
rect 1582 0 1638 400
rect 1950 0 2006 400
rect 2318 0 2374 400
rect 2594 0 2650 400
rect 258 572 366 1604
rect 998 1116 1106 2148
<< via2 >>
rect 940 2202 996 2204
rect 1020 2202 1076 2204
rect 1100 2202 1156 2204
rect 940 2150 978 2202
rect 978 2150 990 2202
rect 990 2150 996 2202
rect 1020 2150 1042 2202
rect 1042 2150 1054 2202
rect 1054 2150 1076 2202
rect 1100 2150 1106 2202
rect 1106 2150 1118 2202
rect 1118 2150 1156 2202
rect 940 2148 996 2150
rect 1020 2148 1076 2150
rect 1100 2148 1156 2150
rect 2340 2202 2396 2204
rect 2420 2202 2476 2204
rect 2500 2202 2556 2204
rect 2340 2150 2378 2202
rect 2378 2150 2390 2202
rect 2390 2150 2396 2202
rect 2420 2150 2442 2202
rect 2442 2150 2454 2202
rect 2454 2150 2476 2202
rect 2500 2150 2506 2202
rect 2506 2150 2518 2202
rect 2518 2150 2556 2202
rect 2340 2148 2396 2150
rect 2420 2148 2476 2150
rect 2500 2148 2556 2150
rect 240 1658 296 1660
rect 320 1658 376 1660
rect 400 1658 456 1660
rect 240 1606 278 1658
rect 278 1606 290 1658
rect 290 1606 296 1658
rect 320 1606 342 1658
rect 342 1606 354 1658
rect 354 1606 376 1658
rect 400 1606 406 1658
rect 406 1606 418 1658
rect 418 1606 456 1658
rect 240 1604 296 1606
rect 320 1604 376 1606
rect 400 1604 456 1606
rect 1640 1658 1696 1660
rect 1720 1658 1776 1660
rect 1800 1658 1856 1660
rect 1640 1606 1678 1658
rect 1678 1606 1690 1658
rect 1690 1606 1696 1658
rect 1720 1606 1742 1658
rect 1742 1606 1754 1658
rect 1754 1606 1776 1658
rect 1800 1606 1806 1658
rect 1806 1606 1818 1658
rect 1818 1606 1856 1658
rect 1640 1604 1696 1606
rect 1720 1604 1776 1606
rect 1800 1604 1856 1606
rect 940 1114 996 1116
rect 1020 1114 1076 1116
rect 1100 1114 1156 1116
rect 940 1062 978 1114
rect 978 1062 990 1114
rect 990 1062 996 1114
rect 1020 1062 1042 1114
rect 1042 1062 1054 1114
rect 1054 1062 1076 1114
rect 1100 1062 1106 1114
rect 1106 1062 1118 1114
rect 1118 1062 1156 1114
rect 940 1060 996 1062
rect 1020 1060 1076 1062
rect 1100 1060 1156 1062
rect 2340 1114 2396 1116
rect 2420 1114 2476 1116
rect 2500 1114 2556 1116
rect 2340 1062 2378 1114
rect 2378 1062 2390 1114
rect 2390 1062 2396 1114
rect 2420 1062 2442 1114
rect 2442 1062 2454 1114
rect 2454 1062 2476 1114
rect 2500 1062 2506 1114
rect 2506 1062 2518 1114
rect 2518 1062 2556 1114
rect 2340 1060 2396 1062
rect 2420 1060 2476 1062
rect 2500 1060 2556 1062
rect 240 570 296 572
rect 320 570 376 572
rect 400 570 456 572
rect 240 518 278 570
rect 278 518 290 570
rect 290 518 296 570
rect 320 518 342 570
rect 342 518 354 570
rect 354 518 376 570
rect 400 518 406 570
rect 406 518 418 570
rect 418 518 456 570
rect 240 516 296 518
rect 320 516 376 518
rect 400 516 456 518
rect 1640 570 1696 572
rect 1720 570 1776 572
rect 1800 570 1856 572
rect 1640 518 1678 570
rect 1678 518 1690 570
rect 1690 518 1696 570
rect 1720 518 1742 570
rect 1742 518 1754 570
rect 1754 518 1776 570
rect 1800 518 1806 570
rect 1806 518 1818 570
rect 1818 518 1856 570
rect 1640 516 1696 518
rect 1720 516 1776 518
rect 1800 516 1856 518
<< metal3 >>
rect 208 496 1888 592
rect 908 1040 2588 1136
rect 208 1584 1888 1680
rect 908 2128 2588 2224
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 276 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 276 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1715205430
transform 1 0 2116 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1715205430
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1715205430
transform 1 0 1932 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[1\]
timestamp 1715205430
transform 1 0 644 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[2\]
timestamp 1715205430
transform 1 0 920 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[3\]
timestamp 1715205430
transform 1 0 1196 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[4\]
timestamp 1715205430
transform 1 0 1472 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[5\]
timestamp 1715205430
transform 1 0 1748 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[6\]
timestamp 1715205430
transform 1 0 2208 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[7\]
timestamp 1715205430
transform 1 0 2484 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 0 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1715205430
transform -1 0 3204 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1715205430
transform 1 0 0 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1715205430
transform -1 0 2760 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1715205430
transform 1 0 0 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1715205430
transform -1 0 3204 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0
timestamp 1715205430
transform -1 0 3204 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1715205430
transform 1 0 2116 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1715205430
transform 1 0 276 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1715205430
transform 1 0 1932 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0
timestamp 1715205430
transform 1 0 2668 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 2024 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_7
timestamp 1715205430
transform -1 0 2928 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_8
timestamp 1715205430
transform 1 0 2836 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_9
timestamp 1715205430
transform 1 0 2024 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_10
timestamp 1715205430
transform 1 0 2836 0 1 1632
box -38 -48 130 592
<< labels >>
flabel metal3 s 208 496 1888 592 0 FreeSans 800 0 0 0 VGND
port 0 nsew ground input
flabel metal3 s 208 1584 1888 1680 0 FreeSans 800 0 0 0 VGND
port 0 nsew ground input
flabel metal3 s 908 1040 2588 1136 0 FreeSans 800 0 0 0 VPWR
port 1 nsew power input
flabel metal3 s 908 2128 2588 2224 0 FreeSans 800 0 0 0 VPWR
port 1 nsew power input
flabel metal2 s 1950 0 2006 400 0 FreeSans 320 90 0 0 gpio_defaults[5]
port 7 nsew signal tristate
flabel metal2 s 2594 0 2650 400 0 FreeSans 320 90 0 0 gpio_defaults[7]
port 9 nsew signal tristate
flabel metal2 s 2318 0 2374 400 0 FreeSans 320 90 0 0 gpio_defaults[6]
port 8 nsew signal tristate
flabel metal2 s 1582 0 1638 400 0 FreeSans 320 90 0 0 gpio_defaults[4]
port 6 nsew signal tristate
flabel metal2 s 1306 0 1362 400 0 FreeSans 320 90 0 0 gpio_defaults[3]
port 5 nsew signal tristate
flabel metal2 s 1030 0 1086 400 0 FreeSans 320 90 0 0 gpio_defaults[2]
port 4 nsew signal tristate
flabel metal2 s 754 0 810 400 0 FreeSans 320 90 0 0 gpio_defaults[1]
port 3 nsew signal tristate
flabel metal2 s 478 0 534 400 0 FreeSans 320 90 0 0 gpio_defaults[0]
port 2 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 3204 2200
<< end >>
